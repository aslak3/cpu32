library IEEE;
use IEEE.STD_LOGIC_1164.all;

package P_CONTROL is
	subtype T_OPCODE is STD_LOGIC_VECTOR (7 downto 0);

	type T_ALU_REG2_MUX_SEL is
		( S_INSTRUCTION_REG2, S_PC );
	type T_ALU_REG3_MUX_SEL is
		( S_INSTRUCTION_REG3, S_INSTRUCTION_QUICK_BYTENYBBLE, S_DATA_IN );
	type T_ALU_OP_MUX_SEL is
		( S_INSTRUCTION_ALU_OP, S_ADD );
	type T_REGS_INPUT_MUX_SEL is
		( S_ALU_RESULT, S_DATA_IN, S_INSTRUCTION_REG2, S_INSTRUCTION_QUICK_WORD );
	type T_REGS_WRITE_INDEX_MUX_SEL is
		( S_INSTRUCTION_REG1, S_STACK_MULTI );
	type T_REGS_READ_REG1_INDEX_MUX_SEL is
		( S_INSTRUCTION_REG1, S_STACK_MULTI );
	type T_PC_INPUT_MUX_SEL is
		( S_ALU_RESULT, S_DATA_IN, S_TEMPORARY_OUTPUT, S_INSTRUCTION_REG1 );
	type T_TEMPORARY_INPUT_MUX_SEL is
		( S_ALU_RESULT, S_DATA_IN );
	type T_ADDRESS_MUX_SEL is
		( S_PC, S_INSTRUCTION_REG2, S_ALU_RESULT, S_TEMPORARY_OUTPUT );
	type T_DATA_OUT_MUX_SEL is
		( S_PC, S_INSTRUCTION_REG1 );

	subtype T_CONDITION is STD_LOGIC_VECTOR (3 downto 0);
end package;
